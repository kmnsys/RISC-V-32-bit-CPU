module InsDec_tb();
    reg [31:0] IR;
    reg [4:0] num ;
    wire MA, MB, MD, RW, MW, MR, PL, JL, JLR, BR;
    wire [3:0] FS;
    wire [2:0] BMC;
    wire [4:0] AA, BA, DA;
    
    
    InsDec UUT(
        .IR(IR),
        .MA(MA), .MB(MB), .MD(MD), .MR(MR),
        .RW(RW), .MW(MW), 
        .PL(PL), .JL(JL), .JLR(JLR), .BR(BR),
        .FS(FS), .BMC(BMC),
        .AA(AA), .BA(BA), .DA(DA)
    );
    
    parameter clk_per = 20;
    
    //rs1:t5-00101
    //rs2:t6-00110
    //rd:t7-00111
    initial begin
    
        //LUI&AUIPC
		#(clk_per);
		IR = 32'b00000000000000000000001110110111;    //lui
		num = 1;
		#(clk_per);
		IR = 32'b00000000000000000000001110010111;    //auipc
		num = 2;
		
		//JUMP&LINK
		#(clk_per);
		IR = 32'b00000000000000000000001111101111;    //jal
		num = 3;
		#(clk_per);
		IR = 32'b00000000000000101000001111100111;    //jlr
		num = 4;
		
		//BRANCHES
		#(clk_per);
		IR = 32'b00000000011000101000000001100011;    //beq
		num = 5;
		#(clk_per);
		IR = 32'b00000000011000101001000001100011;    //bne
		num = 6;
		#(clk_per);
		IR = 32'b00000000011000101100000001100011;    //blt
		num = 7;
		#(clk_per);
		IR = 32'b00000000011000101101000001100011;    //bge
		num = 8;
		#(clk_per);
		IR = 32'b00000000011000101110000001100011;    //bltu
		num = 9;
		#(clk_per);
		IR = 32'b00000000011000101111000001100011;    //bgeu
		num = 10;
		
        //LOADS
		#(clk_per);
		IR = 32'b00000000000000101000001110000011;    //lb 
		num = 11;
		#(clk_per);
		IR = 32'b00000000000000101001001110000011;    //lh 
		num = 12;
		#(clk_per);
		IR = 32'b00000000000000101010001110000011;    //lw 
		num = 13;
		#(clk_per);
		IR = 32'b00000000000000101100001110000011;    //lbu
		num = 14;
		#(clk_per); 
		IR = 32'b00000000000000101101001110000011;    //lhu
		num = 15;
		
		//STORES
		#(clk_per);
		IR = 32'b00000000011000101000000000100011;    //sb
		num = 16;
		#(clk_per);
		IR = 32'b00000000011000101001000000100011;    //sh
		num = 17;
		#(clk_per);
		IR = 32'b00000000011000101010000000100011;    //sw
		num = 18;
        
		//FU IMM
		#(clk_per);
		IR = 32'b00000000000000101000001110010011;    //addi
		num = 19;
		#(clk_per);
		IR = 32'b00000000000000101010001110010011;    //slti
		num = 20;
		#(clk_per);
		IR = 32'b00000000000000101011001110010011;    //stiu
		num = 21;
		#(clk_per);
		IR = 32'b00000000000000101100001110010011;    //xori
		num = 22;
		#(clk_per);
		IR = 32'b00000000000000101110001110010011;    //ori
		num = 23;
		#(clk_per);
		IR = 32'b00000000000000101111001110010011;    //andi
		num = 24;
		#(clk_per);
		IR = 32'b00000000000000101001001110010011;    //slli
		num = 25;
		#(clk_per);
		IR = 32'b00000000000000101101001110010011;    //srli
		num = 26;
		#(clk_per);
		IR = 32'b01000000000000101101001110010011;    //srai
		num = 27;
        
		//FU
		#(clk_per);
		IR = 32'b00000000011000101000001110110011;    //add
		num = 28;
		#(clk_per);
		IR = 32'b01000000011000101000001110110011;    //sub
		num = 29;
		#(clk_per);
		IR = 32'b00000000011000101001001110110011;    //sll
		num = 30;
		#(clk_per);
		IR = 32'b00000000011000101010001110110011;    //slt
		num = 31;
		#(clk_per);
		IR = 32'b00000000011000101011001110110011;    //sltu
		num = 32;
		#(clk_per);
		IR = 32'b00000000011000101100001110110011;    //xor
		num = 33;
		#(clk_per);
		IR = 32'b00000000011000101101001110110011;    //srl
		num = 34;
		#(clk_per);
		IR = 32'b01000000011000101101001110110011;    //sra
		num = 35;
		#(clk_per);
		IR = 32'b00000000011000101110001110110011;    //or
		num = 36;
		#(clk_per);
		IR = 32'b00000000011000101111001110110011;    //and
		num = 37;
		#(clk_per);
		
		$finish;
    
    end
endmodule
